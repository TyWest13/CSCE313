// nios_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nios_system (
		input  wire [3:0]  bcdin_export,   //   bcdin.export
		input  wire        clk_clk,        //     clk.clk
		output wire [7:0]  cout_export,    //    cout.export
		input  wire [1:0]  modes_export,   //   modes.export
		output wire [17:0] pattern_export, // pattern.export
		input  wire        reset_reset_n,  //   reset.reset_n
		output wire [7:0]  seg0_export,    //    seg0.export
		output wire [7:0]  seg1_export,    //    seg1.export
		output wire [7:0]  seg2_export,    //    seg2.export
		output wire [7:0]  seg3_export,    //    seg3.export
		output wire [7:0]  seg4_export,    //    seg4.export
		input  wire        spcont_export   //  spcont.export
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [17:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                      // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [17:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;               // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] mm_interconnect_0_system_modes_s1_readdata;                  // system_modes:readdata -> mm_interconnect_0:system_modes_s1_readdata
	wire   [1:0] mm_interconnect_0_system_modes_s1_address;                   // mm_interconnect_0:system_modes_s1_address -> system_modes:address
	wire         mm_interconnect_0_system_counter_s1_chipselect;              // mm_interconnect_0:system_counter_s1_chipselect -> system_counter:chipselect
	wire  [31:0] mm_interconnect_0_system_counter_s1_readdata;                // system_counter:readdata -> mm_interconnect_0:system_counter_s1_readdata
	wire   [1:0] mm_interconnect_0_system_counter_s1_address;                 // mm_interconnect_0:system_counter_s1_address -> system_counter:address
	wire         mm_interconnect_0_system_counter_s1_write;                   // mm_interconnect_0:system_counter_s1_write -> system_counter:write_n
	wire  [31:0] mm_interconnect_0_system_counter_s1_writedata;               // mm_interconnect_0:system_counter_s1_writedata -> system_counter:writedata
	wire         mm_interconnect_0_random_pattern_s1_chipselect;              // mm_interconnect_0:random_pattern_s1_chipselect -> random_pattern:chipselect
	wire  [31:0] mm_interconnect_0_random_pattern_s1_readdata;                // random_pattern:readdata -> mm_interconnect_0:random_pattern_s1_readdata
	wire   [1:0] mm_interconnect_0_random_pattern_s1_address;                 // mm_interconnect_0:random_pattern_s1_address -> random_pattern:address
	wire         mm_interconnect_0_random_pattern_s1_write;                   // mm_interconnect_0:random_pattern_s1_write -> random_pattern:write_n
	wire  [31:0] mm_interconnect_0_random_pattern_s1_writedata;               // mm_interconnect_0:random_pattern_s1_writedata -> random_pattern:writedata
	wire         mm_interconnect_0_segment0_s1_chipselect;                    // mm_interconnect_0:segment0_s1_chipselect -> segment0:chipselect
	wire  [31:0] mm_interconnect_0_segment0_s1_readdata;                      // segment0:readdata -> mm_interconnect_0:segment0_s1_readdata
	wire   [1:0] mm_interconnect_0_segment0_s1_address;                       // mm_interconnect_0:segment0_s1_address -> segment0:address
	wire         mm_interconnect_0_segment0_s1_write;                         // mm_interconnect_0:segment0_s1_write -> segment0:write_n
	wire  [31:0] mm_interconnect_0_segment0_s1_writedata;                     // mm_interconnect_0:segment0_s1_writedata -> segment0:writedata
	wire         mm_interconnect_0_segment1_s1_chipselect;                    // mm_interconnect_0:segment1_s1_chipselect -> segment1:chipselect
	wire  [31:0] mm_interconnect_0_segment1_s1_readdata;                      // segment1:readdata -> mm_interconnect_0:segment1_s1_readdata
	wire   [1:0] mm_interconnect_0_segment1_s1_address;                       // mm_interconnect_0:segment1_s1_address -> segment1:address
	wire         mm_interconnect_0_segment1_s1_write;                         // mm_interconnect_0:segment1_s1_write -> segment1:write_n
	wire  [31:0] mm_interconnect_0_segment1_s1_writedata;                     // mm_interconnect_0:segment1_s1_writedata -> segment1:writedata
	wire         mm_interconnect_0_segment2_s1_chipselect;                    // mm_interconnect_0:segment2_s1_chipselect -> segment2:chipselect
	wire  [31:0] mm_interconnect_0_segment2_s1_readdata;                      // segment2:readdata -> mm_interconnect_0:segment2_s1_readdata
	wire   [1:0] mm_interconnect_0_segment2_s1_address;                       // mm_interconnect_0:segment2_s1_address -> segment2:address
	wire         mm_interconnect_0_segment2_s1_write;                         // mm_interconnect_0:segment2_s1_write -> segment2:write_n
	wire  [31:0] mm_interconnect_0_segment2_s1_writedata;                     // mm_interconnect_0:segment2_s1_writedata -> segment2:writedata
	wire         mm_interconnect_0_segment3_s1_chipselect;                    // mm_interconnect_0:segment3_s1_chipselect -> segment3:chipselect
	wire  [31:0] mm_interconnect_0_segment3_s1_readdata;                      // segment3:readdata -> mm_interconnect_0:segment3_s1_readdata
	wire   [1:0] mm_interconnect_0_segment3_s1_address;                       // mm_interconnect_0:segment3_s1_address -> segment3:address
	wire         mm_interconnect_0_segment3_s1_write;                         // mm_interconnect_0:segment3_s1_write -> segment3:write_n
	wire  [31:0] mm_interconnect_0_segment3_s1_writedata;                     // mm_interconnect_0:segment3_s1_writedata -> segment3:writedata
	wire         mm_interconnect_0_segment4_s1_chipselect;                    // mm_interconnect_0:segment4_s1_chipselect -> segment4:chipselect
	wire  [31:0] mm_interconnect_0_segment4_s1_readdata;                      // segment4:readdata -> mm_interconnect_0:segment4_s1_readdata
	wire   [1:0] mm_interconnect_0_segment4_s1_address;                       // mm_interconnect_0:segment4_s1_address -> segment4:address
	wire         mm_interconnect_0_segment4_s1_write;                         // mm_interconnect_0:segment4_s1_write -> segment4:write_n
	wire  [31:0] mm_interconnect_0_segment4_s1_writedata;                     // mm_interconnect_0:segment4_s1_writedata -> segment4:writedata
	wire  [31:0] mm_interconnect_0_bcd_input_s1_readdata;                     // bcd_input:readdata -> mm_interconnect_0:bcd_input_s1_readdata
	wire   [1:0] mm_interconnect_0_bcd_input_s1_address;                      // mm_interconnect_0:bcd_input_s1_address -> bcd_input:address
	wire  [31:0] mm_interconnect_0_speed_controller_s1_readdata;              // speed_controller:readdata -> mm_interconnect_0:speed_controller_s1_readdata
	wire   [1:0] mm_interconnect_0_speed_controller_s1_address;               // mm_interconnect_0:speed_controller_s1_address -> speed_controller:address
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [bcd_input:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, random_pattern:reset_n, rst_translator:in_reset, segment0:reset_n, segment1:reset_n, segment2:reset_n, segment3:reset_n, segment4:reset_n, speed_controller:reset_n, system_counter:reset_n, system_modes:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	nios_system_bcd_input bcd_input (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_bcd_input_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_bcd_input_s1_readdata), //                    .readdata
		.in_port  (bcdin_export)                             // external_connection.export
	);

	nios_system_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_system_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	nios_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	nios_system_random_pattern random_pattern (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_random_pattern_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_random_pattern_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_random_pattern_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_random_pattern_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_random_pattern_s1_readdata),   //                    .readdata
		.out_port   (pattern_export)                                  // external_connection.export
	);

	nios_system_segment0 segment0 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_segment0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segment0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segment0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segment0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segment0_s1_readdata),   //                    .readdata
		.out_port   (seg0_export)                               // external_connection.export
	);

	nios_system_segment0 segment1 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_segment1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segment1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segment1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segment1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segment1_s1_readdata),   //                    .readdata
		.out_port   (seg1_export)                               // external_connection.export
	);

	nios_system_segment0 segment2 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_segment2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segment2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segment2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segment2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segment2_s1_readdata),   //                    .readdata
		.out_port   (seg2_export)                               // external_connection.export
	);

	nios_system_segment0 segment3 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_segment3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segment3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segment3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segment3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segment3_s1_readdata),   //                    .readdata
		.out_port   (seg3_export)                               // external_connection.export
	);

	nios_system_segment0 segment4 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_segment4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segment4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segment4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segment4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segment4_s1_readdata),   //                    .readdata
		.out_port   (seg4_export)                               // external_connection.export
	);

	nios_system_speed_controller speed_controller (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_speed_controller_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_speed_controller_s1_readdata), //                    .readdata
		.in_port  (spcont_export)                                   // external_connection.export
	);

	nios_system_segment0 system_counter (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_system_counter_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_system_counter_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_system_counter_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_system_counter_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_system_counter_s1_readdata),   //                    .readdata
		.out_port   (cout_export)                                     // external_connection.export
	);

	nios_system_system_modes system_modes (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_system_modes_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_system_modes_s1_readdata), //                    .readdata
		.in_port  (modes_export)                                // external_connection.export
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_readdatavalid         (nios2_gen2_0_data_master_readdatavalid),                      //                                         .readdatavalid
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.nios2_gen2_0_instruction_master_readdatavalid  (nios2_gen2_0_instruction_master_readdatavalid),               //                                         .readdatavalid
		.bcd_input_s1_address                           (mm_interconnect_0_bcd_input_s1_address),                      //                             bcd_input_s1.address
		.bcd_input_s1_readdata                          (mm_interconnect_0_bcd_input_s1_readdata),                     //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.random_pattern_s1_address                      (mm_interconnect_0_random_pattern_s1_address),                 //                        random_pattern_s1.address
		.random_pattern_s1_write                        (mm_interconnect_0_random_pattern_s1_write),                   //                                         .write
		.random_pattern_s1_readdata                     (mm_interconnect_0_random_pattern_s1_readdata),                //                                         .readdata
		.random_pattern_s1_writedata                    (mm_interconnect_0_random_pattern_s1_writedata),               //                                         .writedata
		.random_pattern_s1_chipselect                   (mm_interconnect_0_random_pattern_s1_chipselect),              //                                         .chipselect
		.segment0_s1_address                            (mm_interconnect_0_segment0_s1_address),                       //                              segment0_s1.address
		.segment0_s1_write                              (mm_interconnect_0_segment0_s1_write),                         //                                         .write
		.segment0_s1_readdata                           (mm_interconnect_0_segment0_s1_readdata),                      //                                         .readdata
		.segment0_s1_writedata                          (mm_interconnect_0_segment0_s1_writedata),                     //                                         .writedata
		.segment0_s1_chipselect                         (mm_interconnect_0_segment0_s1_chipselect),                    //                                         .chipselect
		.segment1_s1_address                            (mm_interconnect_0_segment1_s1_address),                       //                              segment1_s1.address
		.segment1_s1_write                              (mm_interconnect_0_segment1_s1_write),                         //                                         .write
		.segment1_s1_readdata                           (mm_interconnect_0_segment1_s1_readdata),                      //                                         .readdata
		.segment1_s1_writedata                          (mm_interconnect_0_segment1_s1_writedata),                     //                                         .writedata
		.segment1_s1_chipselect                         (mm_interconnect_0_segment1_s1_chipselect),                    //                                         .chipselect
		.segment2_s1_address                            (mm_interconnect_0_segment2_s1_address),                       //                              segment2_s1.address
		.segment2_s1_write                              (mm_interconnect_0_segment2_s1_write),                         //                                         .write
		.segment2_s1_readdata                           (mm_interconnect_0_segment2_s1_readdata),                      //                                         .readdata
		.segment2_s1_writedata                          (mm_interconnect_0_segment2_s1_writedata),                     //                                         .writedata
		.segment2_s1_chipselect                         (mm_interconnect_0_segment2_s1_chipselect),                    //                                         .chipselect
		.segment3_s1_address                            (mm_interconnect_0_segment3_s1_address),                       //                              segment3_s1.address
		.segment3_s1_write                              (mm_interconnect_0_segment3_s1_write),                         //                                         .write
		.segment3_s1_readdata                           (mm_interconnect_0_segment3_s1_readdata),                      //                                         .readdata
		.segment3_s1_writedata                          (mm_interconnect_0_segment3_s1_writedata),                     //                                         .writedata
		.segment3_s1_chipselect                         (mm_interconnect_0_segment3_s1_chipselect),                    //                                         .chipselect
		.segment4_s1_address                            (mm_interconnect_0_segment4_s1_address),                       //                              segment4_s1.address
		.segment4_s1_write                              (mm_interconnect_0_segment4_s1_write),                         //                                         .write
		.segment4_s1_readdata                           (mm_interconnect_0_segment4_s1_readdata),                      //                                         .readdata
		.segment4_s1_writedata                          (mm_interconnect_0_segment4_s1_writedata),                     //                                         .writedata
		.segment4_s1_chipselect                         (mm_interconnect_0_segment4_s1_chipselect),                    //                                         .chipselect
		.speed_controller_s1_address                    (mm_interconnect_0_speed_controller_s1_address),               //                      speed_controller_s1.address
		.speed_controller_s1_readdata                   (mm_interconnect_0_speed_controller_s1_readdata),              //                                         .readdata
		.system_counter_s1_address                      (mm_interconnect_0_system_counter_s1_address),                 //                        system_counter_s1.address
		.system_counter_s1_write                        (mm_interconnect_0_system_counter_s1_write),                   //                                         .write
		.system_counter_s1_readdata                     (mm_interconnect_0_system_counter_s1_readdata),                //                                         .readdata
		.system_counter_s1_writedata                    (mm_interconnect_0_system_counter_s1_writedata),               //                                         .writedata
		.system_counter_s1_chipselect                   (mm_interconnect_0_system_counter_s1_chipselect),              //                                         .chipselect
		.system_modes_s1_address                        (mm_interconnect_0_system_modes_s1_address),                   //                          system_modes_s1.address
		.system_modes_s1_readdata                       (mm_interconnect_0_system_modes_s1_readdata)                   //                                         .readdata
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
